* simulation file template for Hibikino
****
* copy from *.cex here (except .end)

****
vji 3 0 pwl 0ns 0v 100ns 0v 101ns 5v 200ns 5v
vs 1 0 dc 5v
.tran 1ns 200ns
.end
